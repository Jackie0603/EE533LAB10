// 64Width 256Deep

// D_Mem u_DMem (.addra(rdata1_Stg3),.addrb(rdata2_Stg3),.clka(clk),.clkb(clk),
              //.dinb(rdata2_Stg3),.douta(Mem_out_Stg3),.web(WMemEn_Stg3));

module D_Mem(
// a - Read    b - Write
input [7:0] addra, addrb,
input rst,
input clka, clkb,
input [63:0] dinb, // write data
output reg [63:0] douta,
input web

);

reg [63:0] D_bram [255:0];

integer i;
always@(posedge clkb or posedge rst)begin
if(rst) begin
    D_bram[0] <= 64'd4;
    D_bram[1] <= 64'd0;
    D_bram[2] <= 64'd0;
    D_bram[3] <= 64'd0;
    D_bram[4] <= 64'd100;
    D_bram[5] <= 64'd0;
    D_bram[6] <= 64'd0;
    D_bram[7] <= 64'd0;
    D_bram[8] <= 64'd0;
    D_bram[9] <= 64'd0;
    D_bram[10] <= 64'd0;
    D_bram[11] <= 64'd0;
    D_bram[12] <= 64'd0;
    D_bram[13] <= 64'd0;
    D_bram[14] <= 64'd0;
    D_bram[15] <= 64'd0;
    D_bram[16] <= 64'd0;
    D_bram[17] <= 64'd0;
    D_bram[18] <= 64'd0;
    D_bram[19] <= 64'd0;
    D_bram[20] <= 64'd0;
    D_bram[21] <= 64'd0;
    D_bram[22] <= 64'd0;
    D_bram[23] <= 64'd0;
    D_bram[24] <= 64'd0;
    D_bram[25] <= 64'd0;
    D_bram[26] <= 64'd0;
    D_bram[27] <= 64'd0;
    D_bram[28] <= 64'd0;
    D_bram[29] <= 64'd0;
    D_bram[30] <= 64'd0;
    D_bram[31] <= 64'd0;
    D_bram[32] <= 64'd0;
    D_bram[33] <= 64'd0;
    D_bram[34] <= 64'd0;
    D_bram[35] <= 64'd0;
    D_bram[36] <= 64'd0;
    D_bram[37] <= 64'd0;
    D_bram[38] <= 64'd0;
    D_bram[39] <= 64'd0;
    D_bram[40] <= 64'd0;
    D_bram[41] <= 64'd0;
    D_bram[42] <= 64'd0;
    D_bram[43] <= 64'd0;
    D_bram[44] <= 64'd0;
    D_bram[45] <= 64'd0;
    D_bram[46] <= 64'd0;
    D_bram[47] <= 64'd0;
    D_bram[48] <= 64'd0;
    D_bram[49] <= 64'd0;
    D_bram[50] <= 64'd0;
    D_bram[51] <= 64'd0;
    D_bram[52] <= 64'd0;
    D_bram[53] <= 64'd0;
    D_bram[54] <= 64'd0;
    D_bram[55] <= 64'd0;
    D_bram[56] <= 64'd0;
    D_bram[57] <= 64'd0;
    D_bram[58] <= 64'd0;
    D_bram[59] <= 64'd0;
    D_bram[60] <= 64'd0;
    D_bram[61] <= 64'd0;
    D_bram[62] <= 64'd0;
    D_bram[63] <= 64'd0;
    D_bram[64] <= 64'd0;
    D_bram[65] <= 64'd0;
    D_bram[66] <= 64'd0;
    D_bram[67] <= 64'd0;
    D_bram[68] <= 64'd0;
    D_bram[69] <= 64'd0;
    D_bram[70] <= 64'd0;
    D_bram[71] <= 64'd0;
    D_bram[72] <= 64'd0;
    D_bram[73] <= 64'd0;
    D_bram[74] <= 64'd0;
    D_bram[75] <= 64'd0;
    D_bram[76] <= 64'd0;
    D_bram[77] <= 64'd0;
    D_bram[78] <= 64'd0;
    D_bram[79] <= 64'd0;
    D_bram[80] <= 64'd0;
    D_bram[81] <= 64'd0;
    D_bram[82] <= 64'd0;
    D_bram[83] <= 64'd0;
    D_bram[84] <= 64'd0;
    D_bram[85] <= 64'd0;
    D_bram[86] <= 64'd0;
    D_bram[87] <= 64'd0;
    D_bram[88] <= 64'd0;
    D_bram[89] <= 64'd0;
    D_bram[90] <= 64'd0;
    D_bram[91] <= 64'd0;
    D_bram[92] <= 64'd0;
    D_bram[93] <= 64'd0;
    D_bram[94] <= 64'd0;
    D_bram[95] <= 64'd0;
    D_bram[96] <= 64'd0;
    D_bram[97] <= 64'd0;
    D_bram[98] <= 64'd0;
    D_bram[99] <= 64'd0;
    D_bram[100] <= 64'd0;
    D_bram[101] <= 64'd0;
    D_bram[102] <= 64'd0;
    D_bram[103] <= 64'd0;
    D_bram[104] <= 64'd0;
    D_bram[105] <= 64'd0;
    D_bram[106] <= 64'd0;
    D_bram[107] <= 64'd0;
    D_bram[108] <= 64'd0;
    D_bram[109] <= 64'd0;
    D_bram[110] <= 64'd0;
    D_bram[111] <= 64'd0;
    D_bram[112] <= 64'd0;
    D_bram[113] <= 64'd0;
    D_bram[114] <= 64'd0;
    D_bram[115] <= 64'd0;
    D_bram[116] <= 64'd0;
    D_bram[117] <= 64'd0;
    D_bram[118] <= 64'd0;
    D_bram[119] <= 64'd0;
    D_bram[120] <= 64'd0;
    D_bram[121] <= 64'd0;
    D_bram[122] <= 64'd0;
    D_bram[123] <= 64'd0;
    D_bram[124] <= 64'd0;
    D_bram[125] <= 64'd0;
    D_bram[126] <= 64'd0;
    D_bram[127] <= 64'd0;
    D_bram[128] <= 64'd0;
    D_bram[129] <= 64'd0;
    D_bram[130] <= 64'd0;
    D_bram[131] <= 64'd0;
    D_bram[132] <= 64'd0;
    D_bram[133] <= 64'd0;
    D_bram[134] <= 64'd0;
    D_bram[135] <= 64'd0;
    D_bram[136] <= 64'd0;
    D_bram[137] <= 64'd0;
    D_bram[138] <= 64'd0;
    D_bram[139] <= 64'd0;
    D_bram[140] <= 64'd0;
    D_bram[141] <= 64'd0;
    D_bram[142] <= 64'd0;
    D_bram[143] <= 64'd0;
    D_bram[144] <= 64'd0;
    D_bram[145] <= 64'd0;
    D_bram[146] <= 64'd0;
    D_bram[147] <= 64'd0;
    D_bram[148] <= 64'd0;
    D_bram[149] <= 64'd0;
    D_bram[150] <= 64'd0;
    D_bram[151] <= 64'd0;
    D_bram[152] <= 64'd0;
    D_bram[153] <= 64'd0;
    D_bram[154] <= 64'd0;
    D_bram[155] <= 64'd0;
    D_bram[156] <= 64'd0;
    D_bram[157] <= 64'd0;
    D_bram[158] <= 64'd0;
    D_bram[159] <= 64'd0;
    D_bram[160] <= 64'd0;
    D_bram[161] <= 64'd0;
    D_bram[162] <= 64'd0;
    D_bram[163] <= 64'd0;
    D_bram[164] <= 64'd0;
    D_bram[165] <= 64'd0;
    D_bram[166] <= 64'd0;
    D_bram[167] <= 64'd0;
    D_bram[168] <= 64'd0;
    D_bram[169] <= 64'd0;
    D_bram[170] <= 64'd0;
    D_bram[171] <= 64'd0;
    D_bram[172] <= 64'd0;
    D_bram[173] <= 64'd0;
    D_bram[174] <= 64'd0;
    D_bram[175] <= 64'd0;
    D_bram[176] <= 64'd0;
    D_bram[177] <= 64'd0;
    D_bram[178] <= 64'd0;
    D_bram[179] <= 64'd0;
    D_bram[180] <= 64'd0;
    D_bram[181] <= 64'd0;
    D_bram[182] <= 64'd0;
    D_bram[183] <= 64'd0;
    D_bram[184] <= 64'd0;
    D_bram[185] <= 64'd0;
    D_bram[186] <= 64'd0;
    D_bram[187] <= 64'd0;
    D_bram[188] <= 64'd0;
    D_bram[189] <= 64'd0;
    D_bram[190] <= 64'd0;
    D_bram[191] <= 64'd0;
    D_bram[192] <= 64'd0;
    D_bram[193] <= 64'd0;
    D_bram[194] <= 64'd0;
    D_bram[195] <= 64'd0;
    D_bram[196] <= 64'd0;
    D_bram[197] <= 64'd0;
    D_bram[198] <= 64'd0;
    D_bram[199] <= 64'd0;
    D_bram[200] <= 64'd0;
    D_bram[201] <= 64'd0;
    D_bram[202] <= 64'd0;
    D_bram[203] <= 64'd0;
    D_bram[204] <= 64'd0;
    D_bram[205] <= 64'd0;
    D_bram[206] <= 64'd0;
    D_bram[207] <= 64'd0;
    D_bram[208] <= 64'd0;
    D_bram[209] <= 64'd0;
    D_bram[210] <= 64'd0;
    D_bram[211] <= 64'd0;
    D_bram[212] <= 64'd0;
    D_bram[213] <= 64'd0;
    D_bram[214] <= 64'd0;
    D_bram[215] <= 64'd0;
    D_bram[216] <= 64'd0;
    D_bram[217] <= 64'd0;
    D_bram[218] <= 64'd0;
    D_bram[219] <= 64'd0;
    D_bram[220] <= 64'd0;
    D_bram[221] <= 64'd0;
    D_bram[222] <= 64'd0;
    D_bram[223] <= 64'd0;
    D_bram[224] <= 64'd0;
    D_bram[225] <= 64'd0;
    D_bram[226] <= 64'd0;
    D_bram[227] <= 64'd0;
    D_bram[228] <= 64'd0;
    D_bram[229] <= 64'd0;
    D_bram[230] <= 64'd0;
    D_bram[231] <= 64'd0;
    D_bram[232] <= 64'd0;
    D_bram[233] <= 64'd0;
    D_bram[234] <= 64'd0;
    D_bram[235] <= 64'd0;
    D_bram[236] <= 64'd0;
    D_bram[237] <= 64'd0;
    D_bram[238] <= 64'd0;
    D_bram[239] <= 64'd0;
    D_bram[240] <= 64'd0;
    D_bram[241] <= 64'd0;
    D_bram[242] <= 64'd0;
    D_bram[243] <= 64'd0;
    D_bram[244] <= 64'd0;
    D_bram[245] <= 64'd0;
    D_bram[246] <= 64'd0;
    D_bram[247] <= 64'd0;
    D_bram[248] <= 64'd0;
    D_bram[249] <= 64'd0;
    D_bram[250] <= 64'd0;
    D_bram[251] <= 64'd0;
    D_bram[252] <= 64'd0;
    D_bram[253] <= 64'd0;
    D_bram[254] <= 64'd0;
    D_bram[255] <= 64'd0;
end
else if(web) begin
    D_bram[addrb] <= dinb;
end
end

always@(posedge clka or posedge rst)begin
if(rst) 
    douta <= 64'd0;
else
    douta <= D_bram[addra];
end

endmodule